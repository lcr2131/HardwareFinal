//Author: Leonard Robinson
//Modified: December 11, 2012
//Issue queue Draft

class issue_queue;

   q[16] issue queue;

   function allocate ();
   endfunction //
   
   function deallocate ();
   endfunction //
   
   function flush ();
   endfunction //

   function shift ();
   endfunction //   
    
   

endclass // issue_queue

interface top_issue_stage_interface(input bit clk);
